module keyboard(clk,resetn,ps2_clk,ps2_data,ready,code);
    input clk,resetn,ps2_clk,ps2_data;
    output reg ready;
    output reg [7:0] code;

    reg loose;
    reg [9:0] buffer;        // ps2_data bits
    reg [3:0] count;  // count ps2_data bits
    reg [2:0] ps2_clk_sync;

    always @(posedge clk) begin
        ps2_clk_sync <=  {ps2_clk_sync[1:0],ps2_clk};
    end

    wire sampling = ps2_clk_sync[2] & ~ps2_clk_sync[1];

    always @(posedge clk) begin
        if (resetn == 0) begin // reset
            count <= 0;
        end
        else begin
            if (sampling) begin
              if (count == 4'd10) begin
                if ((buffer[0] == 0) &&  // start bit
                    (ps2_data)       &&  // stop bit
                    (^buffer[9:1])) begin      // odd  parity
                    $display("receive %x", buffer[8:1]);
                    code <= buffer[8:1];
                    // add
                    if (buffer[8:0] == 8'hf0) begin
                      loose <= 1'b1;
                      ready <= 1'b0;
                    end else begin
                      if(loose == 1'b0) ready <= 1'b1; 
                      loose <= 1'b0;
                    end
                end
                count <= 0;     // for next
              end else begin
                buffer[count] <= ps2_data;  // store ps2_data
                count <= count + 3'b1;
              end
            end
        end
    end

endmodule