module adder
#(N)
(

);

endmodule