module top(y);
  output [7:0]y;
  assign y = 8'b11111001;
endmodule