module PC (
    input [31:0] inst,
    output [63:0] pc
);
endmodule