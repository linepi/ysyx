module PC (
    input [31:0] inst,
    output [63:0] pc
);
    assign pc = 0;
endmodule