module top(y);
  output [7:0]y;
  assign y = 8'b00000001
endmodule