module control (
    input [31:0] inst,
    output flag
);
    
endmodule