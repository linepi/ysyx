module top(y);
  output [7:0]y;
  assign y = 8'b10000000;
endmodule